library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pkg.all;
use work.op_pkg.all;

entity ctrl is
	port (
		clk         : in std_logic;
		res_n       : in std_logic;
		stall       : in std_logic;

		stall_fetch : out std_logic;
		stall_dec   : out std_logic;
		stall_exec  : out std_logic;
		stall_mem   : out std_logic;
		stall_wb    : out std_logic;

		flush_fetch : out std_logic;
		flush_dec   : out std_logic;
		flush_exec  : out std_logic;
		flush_mem   : out std_logic;
		flush_wb    : out std_logic;

		-- from FWD
		wb_op_exec  : in  wb_op_type;
		exec_op_dec : in  exec_op_type;

		pcsrc_in : in std_logic;
		pcsrc_out : out std_logic
	);
end entity;

architecture rtl of ctrl is
begin
	
--	sync : process(all) is
--		-- Declaration(s)
--	begin
--		if res_n = '0' then
--			
--		elsif rising_edge(clk) then
--			state <= state_next;
--			state_next <= state;
--			
--			if
--			if
--		else;
--	end process;
--	
--	async : process(all) is
--		-- Declaration(s)
--	begin
--		case state is
--		when STATE_FLUSH_BRANCH_HI =>
--			flush_fetch <=  '1';
--			flush_dec <=  '1';
--			flush_exec <=  '1';
--		when STATE_FLUSH_BRANCH_LO =>
--			flush_fetch <=  '0';
--			flush_dec <=  '0';
--			flush_exec <=  '0';
--		when others =>
--			flush_fetch <=  '0';
--			flush_dec <=  '0';
--			flush_exec <=  '0';
--		end case;
--	end process;
	
end architecture;
