library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.mem_pkg.all;
use work.cache_pkg.all;
use work.single_clock_rw_ram_pkg.all;

entity data_st_1w is
	generic (
		SETS_LD  : natural := SETS_LD
	);
	port (
		clk       : in std_logic;

		we        : in std_logic;
		rd        : in std_logic;
		index     : in c_index_type;
		byteena   : in mem_byteena_type;

		data_in   : in mem_data_type;
		data_out  : out mem_data_type
);
end entity;

architecture impl of data_st_1w is
begin

	-- each SRAM instance is used for one byte

	CACHE: for i in 3 downto 0 generate
		CBYTE : single_clock_rw_ram
		generic map (
			ADDR_WIDTH => SETS_LD,
			DATA_WIDTH => 8
		)
		port map (
			clk => clk,
			data_in => data_in(8*(i+1)-1 downto 8*i),
			write_address => index,
			read_address => index,
			we => we and byteena(i),
			data_out => data_out(8*(i+1)-1 downto 8*i)
		);
	end generate;

end architecture;
